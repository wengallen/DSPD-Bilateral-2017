// Output SNR ≥ 40 dB (test pattern provided)
// Latency ~= 70k cycles
// Clock frequency: 100MHz
// Technology: UMC 0.18μm process

// Bilateral Filter
module mul_h(
    i000_n,i001_n,i002_n,i003_n,i004_n,i005_n,i006_n,i007_n,i008_n,i009_n,
    i010_n,i011_n,i012_n,i013_n,i014_n,i015_n,i016_n,i017_n,i018_n,i019_n,
    i020_n,i021_n,i022_n,i023_n,i024_n,i025_n,i026_n,i027_n,i028_n,i029_n,
    i030_n,i031_n,i032_n,i033_n,i034_n,i035_n,i036_n,i037_n,i038_n,i039_n,
    i040_n,i041_n,i042_n,i043_n,i044_n,i045_n,i046_n,i047_n,i048_n,i049_n,
    i050_n,i051_n,i052_n,i053_n,i054_n,i055_n,i056_n,i057_n,i058_n,i059_n,
    i060_n,i061_n,i062_n,i063_n,i064_n,i065_n,i066_n,i067_n,i068_n,i069_n,
    i070_n,i071_n,i072_n,i073_n,i074_n,i075_n,i076_n,i077_n,i078_n,i079_n,
    i080_n,i081_n,i082_n,i083_n,i084_n,i085_n,i086_n,i087_n,i088_n,i089_n,
    i090_n,i091_n,i092_n,i093_n,i094_n,i095_n,i096_n,i097_n,i098_n,i099_n,
    i100_n,i101_n,i102_n,i103_n,i104_n,i105_n,i106_n,i107_n,i108_n,i109_n,
    i110_n,i111_n,i112_n,i113_n,i114_n,i115_n,i116_n,i117_n,i118_n,i119_n,i120_n,
    i000_r,i001_r,i002_r,i003_r,i004_r,i005_r,i006_r,i007_r,i008_r,i009_r,
    i010_r,i011_r,i012_r,i013_r,i014_r,i015_r,i016_r,i017_r,i018_r,i019_r,
    i020_r,i021_r,i022_r,i023_r,i024_r,i025_r,i026_r,i027_r,i028_r,i029_r,
    i030_r,i031_r,i032_r,i033_r,i034_r,i035_r,i036_r,i037_r,i038_r,i039_r,
    i040_r,i041_r,i042_r,i043_r,i044_r,i045_r,i046_r,i047_r,i048_r,i049_r,
    i050_r,i051_r,i052_r,i053_r,i054_r,i055_r,i056_r,i057_r,i058_r,i059_r,
    i060_r,i061_r,i062_r,i063_r,i064_r,i065_r,i066_r,i067_r,i068_r,i069_r,
    i070_r,i071_r,i072_r,i073_r,i074_r,i075_r,i076_r,i077_r,i078_r,i079_r,
    i080_r,i081_r,i082_r,i083_r,i084_r,i085_r,i086_r,i087_r,i088_r,i089_r,
    i090_r,i091_r,i092_r,i093_r,i094_r,i095_r,i096_r,i097_r,i098_r,i099_r,
    i100_r,i101_r,i102_r,i103_r,i104_r,i105_r,i106_r,i107_r,i108_r,i109_r,
    i110_r,i111_r,i112_r,i113_r,i114_r,i115_r,i116_r,i117_r,i118_r,i119_r,i120_r,
    out000,out001,out002,out003,out004,out005,out006,out007,out008,out009,
    out010,out011,out012,out013,out014,out015,out016,out017,out018,out019,
    out020,out021,out022,out023,out024,out025,out026,out027,out028,out029,
    out030,out031,out032,out033,out034,out035,out036,out037,out038,out039,
    out040,out041,out042,out043,out044,out045,out046,out047,out048,out049,
    out050,out051,out052,out053,out054,out055,out056,out057,out058,out059,
    out060,out061,out062,out063,out064,out065,out066,out067,out068,out069,
    out070,out071,out072,out073,out074,out075,out076,out077,out078,out079,
    out080,out081,out082,out083,out084,out085,out086,out087,out088,out089,
    out090,out091,out092,out093,out094,out095,out096,out097,out098,out099,
    out100,out101,out102,out103,out104,out105,out106,out107,out108,out109,
    out110,out111,out112,out113,out114,out115,out116,out117,out118,out119,out120,
    en
);

//==== I/O port ==========================
input  [7:0]  i000_n,i001_n,i002_n,i003_n,i004_n,i005_n,i006_n,i007_n,i008_n,i009_n;
input  [7:0]  i010_n,i011_n,i012_n,i013_n,i014_n,i015_n,i016_n,i017_n,i018_n,i019_n;
input  [7:0]  i020_n,i021_n,i022_n,i023_n,i024_n,i025_n,i026_n,i027_n,i028_n,i029_n;
input  [7:0]  i030_n,i031_n,i032_n,i033_n,i034_n,i035_n,i036_n,i037_n,i038_n,i039_n;
input  [7:0]  i040_n,i041_n,i042_n,i043_n,i044_n,i045_n,i046_n,i047_n,i048_n,i049_n;
input  [7:0]  i050_n,i051_n,i052_n,i053_n,i054_n,i055_n,i056_n,i057_n,i058_n,i059_n;
input  [7:0]  i060_n,i061_n,i062_n,i063_n,i064_n,i065_n,i066_n,i067_n,i068_n,i069_n;
input  [7:0]  i070_n,i071_n,i072_n,i073_n,i074_n,i075_n,i076_n,i077_n,i078_n,i079_n;
input  [7:0]  i080_n,i081_n,i082_n,i083_n,i084_n,i085_n,i086_n,i087_n,i088_n,i089_n;
input  [7:0]  i090_n,i091_n,i092_n,i093_n,i094_n,i095_n,i096_n,i097_n,i098_n,i099_n;
input  [7:0]  i100_n,i101_n,i102_n,i103_n,i104_n,i105_n,i106_n,i107_n,i108_n,i109_n;
input  [7:0]  i110_n,i111_n,i112_n,i113_n,i114_n,i115_n,i116_n,i117_n,i118_n,i119_n,i120_n;

input  [13:0] i000_r,i001_r,i002_r,i003_r,i004_r,i005_r,i006_r,i007_r,i008_r,i009_r;
input  [13:0] i010_r,i011_r,i012_r,i013_r,i014_r,i015_r,i016_r,i017_r,i018_r,i019_r;
input  [13:0] i020_r,i021_r,i022_r,i023_r,i024_r,i025_r,i026_r,i027_r,i028_r,i029_r;
input  [13:0] i030_r,i031_r,i032_r,i033_r,i034_r,i035_r,i036_r,i037_r,i038_r,i039_r;
input  [13:0] i040_r,i041_r,i042_r,i043_r,i044_r,i045_r,i046_r,i047_r,i048_r,i049_r;
input  [13:0] i050_r,i051_r,i052_r,i053_r,i054_r,i055_r,i056_r,i057_r,i058_r,i059_r;
input  [13:0] i060_r,i061_r,i062_r,i063_r,i064_r,i065_r,i066_r,i067_r,i068_r,i069_r;
input  [13:0] i070_r,i071_r,i072_r,i073_r,i074_r,i075_r,i076_r,i077_r,i078_r,i079_r;
input  [13:0] i080_r,i081_r,i082_r,i083_r,i084_r,i085_r,i086_r,i087_r,i088_r,i089_r;
input  [13:0] i090_r,i091_r,i092_r,i093_r,i094_r,i095_r,i096_r,i097_r,i098_r,i099_r;
input  [13:0] i100_r,i101_r,i102_r,i103_r,i104_r,i105_r,i106_r,i107_r,i108_r,i109_r;
input  [13:0] i110_r,i111_r,i112_r,i113_r,i114_r,i115_r,i116_r,i117_r,i118_r,i119_r,i120_r;


output reg [27:0] out000,out001,out002,out003,out004,out005,out006,out007,out008,out009;
output reg [27:0] out010,out011,out012,out013,out014,out015,out016,out017,out018,out019;
output reg [27:0] out020,out021,out022,out023,out024,out025,out026,out027,out028,out029;
output reg [27:0] out030,out031,out032,out033,out034,out035,out036,out037,out038,out039;
output reg [27:0] out040,out041,out042,out043,out044,out045,out046,out047,out048,out049;
output reg [27:0] out050,out051,out052,out053,out054,out055,out056,out057,out058,out059;
output reg [27:0] out060,out061,out062,out063,out064,out065,out066,out067,out068,out069;
output reg [27:0] out070,out071,out072,out073,out074,out075,out076,out077,out078,out079;
output reg [27:0] out080,out081,out082,out083,out084,out085,out086,out087,out088,out089;
output reg [27:0] out090,out091,out092,out093,out094,out095,out096,out097,out098,out099;
output reg [27:0] out100,out101,out102,out103,out104,out105,out106,out107,out108,out109;
output reg [27:0] out110,out111,out112,out113,out114,out115,out116,out117,out118,out119,out120;

input         en;

always@(*) begin
    if(en) begin
        out000 = {i000_n,6'b0} * 14'b0_010000;
        out001 = {i001_n,6'b0} * 14'b0_010000;
        out002 = {i002_n,6'b0} * 14'b0_010000;
        out003 = {i003_n,6'b0} * 14'b0_010000;
        out004 = {i004_n,6'b0} * 14'b0_010000;
        out005 = {i005_n,6'b0} * 14'b0_010000;
        out006 = {i006_n,6'b0} * 14'b0_010000;
        out007 = {i007_n,6'b0} * 14'b0_010000;
        out008 = {i008_n,6'b0} * 14'b0_010000;
        out009 = {i009_n,6'b0} * 14'b0_010000;
        out010 = {i010_n,6'b0} * 14'b0_010000;
        out011 = {i011_n,6'b0} * 14'b0_010000;
        out012 = {i012_n,6'b0} * 14'b0_010000;
        out013 = {i013_n,6'b0} * 14'b0_010000;
        out014 = {i014_n,6'b0} * 14'b0_010000;
        out015 = {i015_n,6'b0} * 14'b0_010000;
        out016 = {i016_n,6'b0} * 14'b0_010000;
        out017 = {i017_n,6'b0} * 14'b0_010000;
        out018 = {i018_n,6'b0} * 14'b0_010000;
        out019 = {i019_n,6'b0} * 14'b0_010000;
        out020 = {i020_n,6'b0} * 14'b0_010000;
        out021 = {i021_n,6'b0} * 14'b0_010000;
        out022 = {i022_n,6'b0} * 14'b0_010000;
        out023 = {i023_n,6'b0} * 14'b0_010000;
        out024 = {i024_n,6'b0} * 14'b0_010000;
        out025 = {i025_n,6'b0} * 14'b0_010000;
        out026 = {i026_n,6'b0} * 14'b0_010000;
        out027 = {i027_n,6'b0} * 14'b0_010000;
        out028 = {i028_n,6'b0} * 14'b0_010000;
        out029 = {i029_n,6'b0} * 14'b0_010000;
        out030 = {i030_n,6'b0} * 14'b0_010000;
        out031 = {i031_n,6'b0} * 14'b0_010000;
        out032 = {i032_n,6'b0} * 14'b0_010000;
        out033 = {i033_n,6'b0} * 14'b0_010000;
        out034 = {i034_n,6'b0} * 14'b0_010000;
        out035 = {i035_n,6'b0} * 14'b0_010000;
        out036 = {i036_n,6'b0} * 14'b0_010000;
        out037 = {i037_n,6'b0} * 14'b0_010000;
        out038 = {i038_n,6'b0} * 14'b0_010000;
        out039 = {i039_n,6'b0} * 14'b0_010000;
        out040 = {i040_n,6'b0} * 14'b0_010000;
        out041 = {i041_n,6'b0} * 14'b0_010000;
        out042 = {i042_n,6'b0} * 14'b0_010000;
        out043 = {i043_n,6'b0} * 14'b0_010000;
        out044 = {i044_n,6'b0} * 14'b0_010000;
        out045 = {i045_n,6'b0} * 14'b0_010000;
        out046 = {i046_n,6'b0} * 14'b0_010000;
        out047 = {i047_n,6'b0} * 14'b0_010000;
        out048 = {i048_n,6'b0} * 14'b0_010000;
        out049 = {i049_n,6'b0} * 14'b0_010000;
        out050 = {i050_n,6'b0} * 14'b0_010000;
        out051 = {i051_n,6'b0} * 14'b0_010000;
        out052 = {i052_n,6'b0} * 14'b0_010000;
        out053 = {i053_n,6'b0} * 14'b0_010000;
        out054 = {i054_n,6'b0} * 14'b0_010000;
        out055 = {i055_n,6'b0} * 14'b0_010000;
        out056 = {i056_n,6'b0} * 14'b0_010000;
        out057 = {i057_n,6'b0} * 14'b0_010000;
        out058 = {i058_n,6'b0} * 14'b0_010000;
        out059 = {i059_n,6'b0} * 14'b0_010000;
        out060 = {i060_n,6'b0} * 14'b1_010000;
        out061 = {i061_n,6'b0} * 14'b0_010000;
        out062 = {i062_n,6'b0} * 14'b0_010000;
        out063 = {i063_n,6'b0} * 14'b0_010000;
        out064 = {i064_n,6'b0} * 14'b0_010000;
        out065 = {i065_n,6'b0} * 14'b0_010000;
        out066 = {i066_n,6'b0} * 14'b0_010000;
        out067 = {i067_n,6'b0} * 14'b0_010000;
        out068 = {i068_n,6'b0} * 14'b0_010000;
        out069 = {i069_n,6'b0} * 14'b0_010000;
        out070 = {i070_n,6'b0} * 14'b0_010000;
        out071 = {i071_n,6'b0} * 14'b0_010000;
        out072 = {i072_n,6'b0} * 14'b0_010000;
        out073 = {i073_n,6'b0} * 14'b0_010000;
        out074 = {i074_n,6'b0} * 14'b0_010000;
        out075 = {i075_n,6'b0} * 14'b0_010000;
        out076 = {i076_n,6'b0} * 14'b0_010000;
        out077 = {i077_n,6'b0} * 14'b0_010000;
        out078 = {i078_n,6'b0} * 14'b0_010000;
        out079 = {i079_n,6'b0} * 14'b0_010000;
        out080 = {i080_n,6'b0} * 14'b0_010000;
        out081 = {i081_n,6'b0} * 14'b0_010000;
        out082 = {i082_n,6'b0} * 14'b0_010000;
        out083 = {i083_n,6'b0} * 14'b0_010000;
        out084 = {i084_n,6'b0} * 14'b0_010000;
        out085 = {i085_n,6'b0} * 14'b0_010000;
        out086 = {i086_n,6'b0} * 14'b0_010000;
        out087 = {i087_n,6'b0} * 14'b0_010000;
        out088 = {i088_n,6'b0} * 14'b0_010000;
        out089 = {i089_n,6'b0} * 14'b0_010000;
        out090 = {i090_n,6'b0} * 14'b0_010000;
        out091 = {i091_n,6'b0} * 14'b0_010000;
        out092 = {i092_n,6'b0} * 14'b0_010000;
        out093 = {i093_n,6'b0} * 14'b0_010000;
        out094 = {i094_n,6'b0} * 14'b0_010000;
        out095 = {i095_n,6'b0} * 14'b0_010000;
        out096 = {i096_n,6'b0} * 14'b0_010000;
        out097 = {i097_n,6'b0} * 14'b0_010000;
        out098 = {i098_n,6'b0} * 14'b0_010000;
        out099 = {i099_n,6'b0} * 14'b0_010000;
        out100 = {i100_n,6'b0} * 14'b0_010000;
        out101 = {i101_n,6'b0} * 14'b0_010000;
        out102 = {i102_n,6'b0} * 14'b0_010000;
        out103 = {i103_n,6'b0} * 14'b0_010000;
        out104 = {i104_n,6'b0} * 14'b0_010000;
        out105 = {i105_n,6'b0} * 14'b0_010000;
        out106 = {i106_n,6'b0} * 14'b0_010000;
        out107 = {i107_n,6'b0} * 14'b0_010000;
        out108 = {i108_n,6'b0} * 14'b0_010000;
        out109 = {i109_n,6'b0} * 14'b0_010000;
        out110 = {i110_n,6'b0} * 14'b0_010000;
        out111 = {i111_n,6'b0} * 14'b0_010000;
        out112 = {i112_n,6'b0} * 14'b0_010000;
        out113 = {i113_n,6'b0} * 14'b0_010000;
        out114 = {i114_n,6'b0} * 14'b0_010000;
        out115 = {i115_n,6'b0} * 14'b0_010000;
        out116 = {i116_n,6'b0} * 14'b0_010000;
        out117 = {i117_n,6'b0} * 14'b0_010000;
        out118 = {i118_n,6'b0} * 14'b0_010000;
        out119 = {i119_n,6'b0} * 14'b0_010000;
        out120 = {i120_n,6'b0} * 14'b0_010000;
    end
    else begin
        out000 = {{8'b0,i000_r},6'b0};
        out001 = {{8'b0,i001_r},6'b0};
        out002 = {{8'b0,i002_r},6'b0};
        out003 = {{8'b0,i003_r},6'b0};
        out004 = {{8'b0,i004_r},6'b0};
        out005 = {{8'b0,i005_r},6'b0};
        out006 = {{8'b0,i006_r},6'b0};
        out007 = {{8'b0,i007_r},6'b0};
        out008 = {{8'b0,i008_r},6'b0};
        out009 = {{8'b0,i009_r},6'b0};
        out010 = {{8'b0,i010_r},6'b0};
        out011 = {{8'b0,i011_r},6'b0};
        out012 = {{8'b0,i012_r},6'b0};
        out013 = {{8'b0,i013_r},6'b0};
        out014 = {{8'b0,i014_r},6'b0};
        out015 = {{8'b0,i015_r},6'b0};
        out016 = {{8'b0,i016_r},6'b0};
        out017 = {{8'b0,i017_r},6'b0};
        out018 = {{8'b0,i018_r},6'b0};
        out019 = {{8'b0,i019_r},6'b0};
        out020 = {{8'b0,i020_r},6'b0};
        out021 = {{8'b0,i021_r},6'b0};
        out022 = {{8'b0,i022_r},6'b0};
        out023 = {{8'b0,i023_r},6'b0};
        out024 = {{8'b0,i024_r},6'b0};
        out025 = {{8'b0,i025_r},6'b0};
        out026 = {{8'b0,i026_r},6'b0};
        out027 = {{8'b0,i027_r},6'b0};
        out028 = {{8'b0,i028_r},6'b0};
        out029 = {{8'b0,i029_r},6'b0};
        out030 = {{8'b0,i030_r},6'b0};
        out031 = {{8'b0,i031_r},6'b0};
        out032 = {{8'b0,i032_r},6'b0};
        out033 = {{8'b0,i033_r},6'b0};
        out034 = {{8'b0,i034_r},6'b0};
        out035 = {{8'b0,i035_r},6'b0};
        out036 = {{8'b0,i036_r},6'b0};
        out037 = {{8'b0,i037_r},6'b0};
        out038 = {{8'b0,i038_r},6'b0};
        out039 = {{8'b0,i039_r},6'b0};
        out040 = {{8'b0,i040_r},6'b0};
        out041 = {{8'b0,i041_r},6'b0};
        out042 = {{8'b0,i042_r},6'b0};
        out043 = {{8'b0,i043_r},6'b0};
        out044 = {{8'b0,i044_r},6'b0};
        out045 = {{8'b0,i045_r},6'b0};
        out046 = {{8'b0,i046_r},6'b0};
        out047 = {{8'b0,i047_r},6'b0};
        out048 = {{8'b0,i048_r},6'b0};
        out049 = {{8'b0,i049_r},6'b0};
        out050 = {{8'b0,i050_r},6'b0};
        out051 = {{8'b0,i051_r},6'b0};
        out052 = {{8'b0,i052_r},6'b0};
        out053 = {{8'b0,i053_r},6'b0};
        out054 = {{8'b0,i054_r},6'b0};
        out055 = {{8'b0,i055_r},6'b0};
        out056 = {{8'b0,i056_r},6'b0};
        out057 = {{8'b0,i057_r},6'b0};
        out058 = {{8'b0,i058_r},6'b0};
        out059 = {{8'b0,i059_r},6'b0};
        out060 = {{8'b0,i060_r},6'b0};
        out061 = {{8'b0,i061_r},6'b0};
        out062 = {{8'b0,i062_r},6'b0};
        out063 = {{8'b0,i063_r},6'b0};
        out064 = {{8'b0,i064_r},6'b0};
        out065 = {{8'b0,i065_r},6'b0};
        out066 = {{8'b0,i066_r},6'b0};
        out067 = {{8'b0,i067_r},6'b0};
        out068 = {{8'b0,i068_r},6'b0};
        out069 = {{8'b0,i069_r},6'b0};
        out070 = {{8'b0,i070_r},6'b0};
        out071 = {{8'b0,i071_r},6'b0};
        out072 = {{8'b0,i072_r},6'b0};
        out073 = {{8'b0,i073_r},6'b0};
        out074 = {{8'b0,i074_r},6'b0};
        out075 = {{8'b0,i075_r},6'b0};
        out076 = {{8'b0,i076_r},6'b0};
        out077 = {{8'b0,i077_r},6'b0};
        out078 = {{8'b0,i078_r},6'b0};
        out079 = {{8'b0,i079_r},6'b0};
        out080 = {{8'b0,i080_r},6'b0};
        out081 = {{8'b0,i081_r},6'b0};
        out082 = {{8'b0,i082_r},6'b0};
        out083 = {{8'b0,i083_r},6'b0};
        out084 = {{8'b0,i084_r},6'b0};
        out085 = {{8'b0,i085_r},6'b0};
        out086 = {{8'b0,i086_r},6'b0};
        out087 = {{8'b0,i087_r},6'b0};
        out088 = {{8'b0,i088_r},6'b0};
        out089 = {{8'b0,i089_r},6'b0};
        out090 = {{8'b0,i090_r},6'b0};
        out091 = {{8'b0,i091_r},6'b0};
        out092 = {{8'b0,i092_r},6'b0};
        out093 = {{8'b0,i093_r},6'b0};
        out094 = {{8'b0,i094_r},6'b0};
        out095 = {{8'b0,i095_r},6'b0};
        out096 = {{8'b0,i096_r},6'b0};
        out097 = {{8'b0,i097_r},6'b0};
        out098 = {{8'b0,i098_r},6'b0};
        out099 = {{8'b0,i099_r},6'b0};
        out100 = {{8'b0,i100_r},6'b0};
        out101 = {{8'b0,i101_r},6'b0};
        out102 = {{8'b0,i102_r},6'b0};
        out103 = {{8'b0,i103_r},6'b0};
        out104 = {{8'b0,i104_r},6'b0};
        out105 = {{8'b0,i105_r},6'b0};
        out106 = {{8'b0,i106_r},6'b0};
        out107 = {{8'b0,i107_r},6'b0};
        out108 = {{8'b0,i108_r},6'b0};
        out109 = {{8'b0,i109_r},6'b0};
        out110 = {{8'b0,i110_r},6'b0};
        out111 = {{8'b0,i111_r},6'b0};
        out112 = {{8'b0,i112_r},6'b0};
        out113 = {{8'b0,i113_r},6'b0};
        out114 = {{8'b0,i114_r},6'b0};
        out115 = {{8'b0,i115_r},6'b0};
        out116 = {{8'b0,i116_r},6'b0};
        out117 = {{8'b0,i117_r},6'b0};
        out118 = {{8'b0,i118_r},6'b0};
        out119 = {{8'b0,i119_r},6'b0};
        out120 = {{8'b0,i120_r},6'b0};
    end
end

endmodule